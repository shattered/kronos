library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_textio.all;
use std.textio.all;
use work.uCmdBits.all;
use work.Kronos_Types.all;

entity Microcode is
    port (
        clock   : in std_logic;
        en      : in std_logic;
        addr    : in std_logic_vector(10 downto 0);
	data	: out std_logic_vector(ucmd_bits));
end Microcode;

architecture Behavioral of Microcode is
begin

    process (clock)
        type rom_type is array (0 to 2047) of std_logic_vector (ucmd_bits);
        constant rom : rom_type :=(
            -- microcode start
            "0000000000001111000000000111111111111111",
            "0000000000001001000000000111111111111111",
            "0000000000001111000000000111111111111111",
            "0000000000001111000000000111111111111111",
            "0000000111101000100000000111111111111111",
            "0000000000000001100000000010101010111111",
            "0000000111001001000000000111111111111111",
            "0000000111101000100000000111111111111111",
            "0000000010000001100000000010101111111111",
            "0000000010100001100000000010111111111111",
            "0000000011000001100000000011001111111111",
            "0000000000000001100000000011011111111111",
            "0000000101100001100000000100011111111111",
            "0000000011100001100000000011101111111111",
            "0000000110000001100000000011111111111111",
            "0000000000000001100000000100101111111111",
            "0000000000000001100000000101100111101011",
            "0000000000000001100000111101101111101010",
            "0000000101100001100000101101101111101010",
            "0000111100000011000000000111111111111111",
            "0001000000011011100000000101101111110100",
            "0000000000010101100000000101101111110100",
            "0000000000011011100000000101101111110100",
            "0000000000010101100000000101101111110100",
            "0000000010001111100000000101101111110100",
            "0000000001000001100000000101101111110100",
            "0000000110010000100000000000011111101011",
            "0000000001000001100000000101101111110100",
            "0000000010001101100000000101101111110100",
            "0000000001000001100000000101101111110100",
            "0000000110010000100000000000011111101111",
            "0000000001000001100000000101101111110100",
            "0000000010100001100000000101101111110100",
            "0000000010000111100000000101101111110100",
            "0000000001000001100000000101101111110100",
            "0000000110010000100000000000011111110010",
            "0000000001000001100000000101101111110100",
            "0000000001011011100000000101101111110100",
            "0000000001111101100000000101101111110100",
            "0000000001000001100000000101101111110100",
            "0000000000000001100001110000011001001111",
            "0000000000000001100000000000011010100001",
            "0000000110010000100000000111111111111111",
            "0000000000011011100000000101101111110100",
            "0000000000010101100000000101101111110100",
            "0000000110100110100000000111111111111111",
            "0000000000000001100000000010001111111111",
            "0000000000000001100000000101100101001000",
            "0000000000011011100000000101101111110100",
            "0000000000010101100000000101101111110100",
            "0000000110010000100000000000011111101000",
            "0000000001111011100000000101101111110100",
            "0000000000000001100000000000011010101000",
            "0000000110010000100000000111111111111111",
            "0000000001110011000000000111111111111111",
            "0000000010100001100000000101101111110100",
            "0000000010001101100000000101101111110100",
            "0000000001000001100000000101101111110100",
            "0000000000000001100000000010011111111111",
            "0000000000000001100000000010101111111111",
            "0000000000000001100000000000011010110100",
            "0000000011010001101000111111111111100001",
            "0000000010001011000000000111111111111111",
            "0000000101000010100000000111111111111111",
            "0000000011010001100000000101101111110100",
            "0000000000000001100000000010001111111111",
            "0000000000011011100000000101101111110100",
            "0000000000010101100000000101101111110100",
            "0000000001100001000000000111111111111111",
            "0000000011101111101000111111111111100001",
            "0000000010011001000000000111111111111111",
            "0000000101110100100000000111111111111111",
            "0000000000000001100000110000010000110100",
            "0000000000000001100010000101100100100001",
            "0000000001100001100000000101101111110100",
            "0000000001110101000000000111111111111111",
            "0000000011100101101000111111111111100001",
            "0000000010101011000000000111111111111111",
            "0000000101110100100000000111111111111111",
            "0000000000000001100000110000010000110100",
            "0000000000000001100010000000011010100001",
            "0000000000100001100011110000011111100001",
            "0000000000001001100000000000101111111111",
            "0000000110010010100000000111111111111111",
            "0000000001110101000000000111111111111111",
            "0000000000011011101000111111111111100001",
            "0000000010110111000100000111111111101010",
            "0000000010110011000000000111111111111111",
            "0000000000000001100000000101100100101000",
            "0000000000000011100000110010001111101000",
            "0000000001100001000000000111111111111111",
            "0000000001011111101000111111111111100001",
            "0000000011001011000000000111111111111111",
            "0000000000000001100000000101100000110100",
            "0000000000000001100100000111111111101010",
            "0000000011000011000000000111111111111111",
            "0000000011000101000000000010001111101001",
            "0000000000000001100000000010001010101000",
            "0000000000011011100000000101101111110100",
            "0000000000010101100000000101101111110100",
            "0000000001100001000000000111111111111111",
            "0000000001100001101100111000101111100001",
            "0000000011011011000000000111111111111111",
            "0000000001110011101100111111110000111111",
            "0000000011011011000000000111111111111111",
            "0000000000000001100000000101100000110100",
            "0000000000000011100000110010101111101010",
            "0000000000001001100011111010011111101001",
            "0000000001111001000000100010010001001001",
            "0000000011000011101100111000101111100001",
            "0000000011100111000000000111111111111111",
            "0000000011001101101100111111110000111111",
            "0000000011100111000000000111111111111111",
            "0000000000010101100000110000101111100010",
            "0000000011010011000000000111111111111111",
            "0000000011001111101000111111111111100001",
            "0000000011111011000000000111111111111111",
            "0000000000000001100000000101100000110100",
            "0000000000000001100100000111111111101010",
            "0000000011110011000000000111111111111111",
            "0000000011110101000000000010101111101001",
            "0000000000000001100000000010101010101010",
            "0000000000011011100000000101101111110100",
            "0000000000010101100000000101101111110100",
            "0000000111001001000000000111111111111111",
            "0000000011011001101000111111111111100001",
            "0000000100001111000000000111111111111111",
            "0000000000000001100100000111111111101010",
            "0000000100001011000000000111111111111111",
            "0000000000000001100000000101100000110100",
            "0000000000000001100000000010001111101001",
            "0000000000000001100000000010011111111111",
            "0000000000000001100000000010101111111111",
            "0000000100011100100000000111111111111111",
            "0000000001111001000000000111111111111111",
            "0000000000010101101000111111111111100001",
            "0000000100010101000000000111111111111111",
            "0000000001111001000000000111111111111111",
            "0000000000000001100000000101111111111111",
            "0000000001111111100000000000101111111111",
            "0000000110001000100000000111111111111111",
            "0000000001100001000000000111111111111111",
            "0000000000000001100000000000111111111111",
            "0000000000000001100000000000011010110100",
            "0000000001100001101100111000101111100001",
            "0000000100101101000000000111111111111111",
            "0000000001110011101100111111110000111111",
            "0000000100101101000000000111111111111111",
            "0000000000001001100011111000111111100011",
            "0000000100011111000000100000110001000011",
            "0000000011000011101100111000101111100001",
            "0000000100111001000000000111111111111111",
            "0000000011001101101100111111110000111111",
            "0000000100111001000000000111111111111111",
            "0000000000010101100000110000101111100010",
            "0000000100101001000000000111111111111111",
            "0000000000011011101000111111111111100001",
            "0000000100010101000000000111111111111111",
            "0000000000000001100000000101100001101000",
            "0000000000000011100000110010001111101000",
            "0000000000000000000000000111111111111111",
            "0000000000010001100000000001011111111111",
            "0000000000000001100000000000111111111111",
            "0000000000000001100010010101100010110100",
            "0000000000000001100010011101100001110100",
            "0000000000000001100010100101100001110100",
            "0000000000000001100010101101100001110100",
            "0000000010000001100010110101101111110100",
            "0000000001000001100010111101101111110100",
            "0000000000000001100010111000011010110100",
            "0000000100000001101000011111111111100001",
            "0000000101010011000000000111111111111111",
            "0000000000010001100100011111111111100001",
            "0000000101010011000000000111111111111111",
            "0000000100000001100000000001001111111111",
            "0000000000000001100010000000011010110100",
            "0000000000000001100010000000101010110100",
            "0000000000100001100011110000101111100010",
            "0000000000000001100000100000010001000001",
            "0000000000000001100000000101100000100011",
            "0000000000000011100000110000111111100011",
            "0000000000000011101000111001001111100100",
            "0000000101011111000000000111111111111111",
            "0000000000000011101000111001011111100101",
            "0000000101010011000000000111111111111111",
            "0000000000000000000000000111111111111111",
            "0000000000000001100000000000101010110100",
            "0000000001100001101100111000011111100010",
            "0000000100010101000000000111111111111111",
            "0000000001110101101100111111111111100010",
            "0000001010001101000000000111111111111111",
            "0000000011000011101100111111111111100010",
            "0000000100010101000000000111111111111111",
            "0000000011001111110000111111111111100010",
            "0000000100010101000000000111111111111111",
            "0000000010101110000000111000011111100010",
            "0000000000000001100000000101100001010100",
            "0000000000010001100011110000011111100001",
            "0000000000000101100000000000101111111111",
            "0000000110010011000000000111111111111111",
            "0000000000010001100000000000101111111111",
            "0000000000001001100011111000011111100001",
            "0000000000011111100000011000111111100001",
            "0000000000010101101100111111111111100011",
            "0000000110011101000000000111111111111111",
            "0000000000001111100000110000111111100011",
            "0000000001100001100000110000111111100011",
            "0000000000000001100000000101100001110100",
            "0000000000000011101000111000101111100010",
            "0000000110010011000000000111111111111111",
            "0000000000000000000000000111111111111111",
            "0000000000000001100000010100011111111111",
            "0000000110110100100000000111111111111111",
            "0000000000000001100000000101100101101010",
            "0000000000000001100000001101100110001010",
            "0000000000000001100000010101101001001010",
            "0000000000000001100000011101100110101010",
            "0000000000000000000000100101100111001010",
            "0000000000000001110100000000011111111111",
            "0000000110111101000000000111111111111111",
            "0000000000000001100000000101100000101110",
            "0000000000000010000000110011101111101110",
            "0000000000000011100000000000101111111111",
            "0000000000000001100000000101101000001110",
            "0000000000000001110100110011100001001110",
            "0000000110111111000000110000010001000001",
            "0000000000000001100000000101100000101110",
            "0000000000000010000000110011101111101110",
            "0000000000000001100000011011011010101010",
            "0000000000000001100000101000011010101010",
            "0000000000000001100000000010111010101010",
            "0000000000000001100000000011111010101011",
            "0000000000000001100000010100101010101010",
            "0000000000100001100000111100011111100001",
            "0000000000000001100000001011001010101010",
            "0000000000000001100000100011101010101010",
            "0000000000000011100000111011101111101110",
            "0000000000000001100000000000011010101110",
            "0000000000000001100100000111111111100001",
            "0000001010001101000000000111111111111111",
            "0000000000000011100000111011101111101110",
            "0000000000000011101000111000011111100001",
            "0000000111100001000000000100001010101110",
            "0000000000000000000000000111111111111111",
            "0000000000000001100000000110011111111111",
            "0000000000000001100000000000011111111111",
            "0000000000000011100000000000111111111111",
            "0000000000011001100011111000101111100011",
            "0000000000010011100011111000111111100011",
            "0000000000000001100000000110001111100001",
            "0000000000000011101000111000111111100011",
            "0000000111110011000000110000010001000001",
            "0000000000000001100000000000011111111111",
            "0000000000000011100000000000111111111111",
            "0000000000001101100011111000111111100011",
            "0000000000001111100000100001001111100001",
            "0000000000000001100000000110000010000001",
            "0000000000000011101000111000111111100011",
            "0000000111111111000000110000010001000001",
            "0000000000000111100000100000011111110100",
            "0000000000000001100000000110000000110100",
            "0000000000000000000000000111111111111111",
            "0000000000000111100000000000011111111111",
            "0000001000101001000000000111111111111111",
            "0000000000001111100000000000011111111111",
            "0000001000101001000000000111111111111111",
            "0000000010000011100000000000011111111111",
            "0000001000101001000000000111111111111111",
            "0000000010010011100000000000011111111111",
            "0000001000101001000000000111111111111111",
            "0000000000000001100000000100001111100011",
            "0000000000000001100000000100001111100010",
            "0000000010010101100000000000011111111111",
            "0000001000101001000000000111111111111111",
            "0000001000101010100000000111111111111111",
            "0000111100000011000000000111111111111111",
            "0000000000000001100000000101111111111111",
            "0000000000000001100000110101100000101010",
            "0000000010000001110000111111111111100001",
            "0000001001000101000000000111111111111111",
            "0000000000111111110000111111111111100001",
            "0000001000111111000100000111111111100001",
            "0000001010001101000000000111111111111111",
            "0000000000000011100011111000100000111111",
            "0000000000000001100100011111110110100010",
            "0000001001001001000000000111111111111111",
            "0000001001011111000000000111111111111111",
            "0000000000000011100100011111111111101101",
            "0000001001001001000000000111111111111111",
            "0000001001011111000000000111111111111111",
            "0000000000000001101100110111110110101101",
            "0000001001011101000000000111111111111111",
            "0000000010000011100100101111111111100001",
            "0000001010001101000000000111111111111111",
            "0000000010000101100100101111111111100001",
            "0000001010001101000000000111111111111111",
            "0000000010000111100100101111111111100001",
            "0000001010001101000000000111111111111111",
            "0000000000000001100000000101111111111111",
            "0000000010101001100000000000101111111111",
            "0000000110001000100000000111111111111111",
            "0000111100000011000000000111111111111111",
            "0000000001111111100000000000011111111111",
            "0000000000000001100000110001010000100001",
            "0000000000000001100000001001001010100101",
            "0000001011111111000000000111111111111111",
            "0000000000000001100000000000011111111101",
            "0000000000000011100100011111111111100001",
            "0000001001101111000000000111111111111111",
            "0000000010011001100000000000011111111111",
            "0000001000101001000000000111111111111111",
            "0000000000000101100100011111111111100001",
            "0000001001110111000000000111111111111111",
            "0000000000000111100000000000011111111111",
            "0000001000101001000000000111111111111111",
            "0000000000001001100100011111111111100001",
            "0000001001111111000000000111111111111111",
            "0000000010000001100000000000011111111111",
            "0000001000101001000000000111111111111111",
            "0000000010001011100000000000011111111111",
            "0000001000101001000000000111111111111111",
            "0000000001101111000000000101111111111111",
            "0000111100000011000000000111111111111111",
            "0000001010001101000000000111111001111111",
            "0000000000000001100000000111111111111111",
            "0000000000000001100000000111111111111111",
            "0000000000000000000000000111111111111111",
            "0000001010001101000010000100001001100001",
            "0000000000000001100010000000011001100001",
            "0000000000000001100010000000011001100001",
            "0000001010001101000010000100001001100001",
            "0000000000000011100000111000011111100001",
            "0000000000000001100000000000011010100001",
            "0000000000000001100000000000011010100001",
            "0000000000000001100000110100001001100001",
            "0000000000000000000000000111111111111111",
            "0000001010100101000000000111111111111111",
            "0000001010000111000000000111111001111111",
            "0000000000000001100010111000011001111111",
            "0000000000000001100010000000011001100001",
            "0000001010001001000000110100100000110010",
            "0000111000110111000000000111111111111111",
            "0000001010001101000000000111111001111111",
            "0000001010110011000000000111111111111111",
            "0000001010000111000000000111111001111111",
            "0000000000000001100010111000011001111111",
            "0000000000000001100010000000011001100001",
            "0000001010001001000000111100100000110010",
            "0000111000111111000000000111111111111111",
            "0000001010001101000000000111111001111111",
            "0000000000000000000000000100001010100001",
            "0000000000000000000000000100001010100001",
            "0000000000000011100000111000011111100001",
            "0000000000000001100000000000011010100001",
            "0000000000000001100000000000011010100001",
            "0000000000000001100000110000011001100001",
            "0000000000000000000000000100001010100001",
            "0000000000000000000000000100001010100001",
            "0000000000000000000000000101101000000001",
            "0000000000000000000000000101101000000001",
            "0000000000000011100000111000011111100001",
            "0000000000000001100000000000011010100001",
            "0000000000000001100000000000011010100001",
            "0000000000000001100000110000011001100001",
            "0000000000000000000000000101101000000001",
            "0000000000000001100000110000011001110000",
            "0000000000000000000000000101100001000001",
            "0000000000000001100000000000011010100001",
            "0000000000000000000001111100001111100001",
            "0000000000000000000000000100001010100001",
            "0000000000000001100001110000011000010000",
            "0000000000000001100000000001001010100001",
            "0000000000000001100010000001000001100100",
            "0000000000000000000000000101100010000001",
            "0000000000000001100000110000011000010000",
            "0000000000000000000000000101100001000001",
            "0000000000000001100000000111111111111111",
            "0000000000000001100000000111111111111111",
            "0000000000000001100000000111111111111111",
            "0000000000000001100000000111111111111111",
            "0000000000000001100000000111111111111111",
            "0000000000000000000000000111111111111111",
            "0000000000000001100000000001001111110000",
            "0000000000000001100000000001011010100101",
            "0000000110100110100000000111111111111111",
            "0000000000000001100000000101100101000100",
            "0000000000000001100000000000111111111111",
            "0000000000000001100000001101100101000011",
            "0000000000000001100000000101100010100011",
            "0000000111001001000000000010101111100101",
            "0000000000000001100000000100001010100001",
            "0000000000000000000000000101101111100001",
            "0000000000000011100000111100101111110010",
            "0000001010001011000000000111111111111111",
            "0000001100101101011000000000011111110000",
            "0000001100100011000000000111111111111111",
            "0000000000000001100000111000010000111111",
            "0000000000000001100000111000100001011111",
            "0000000000000001100001010000110001000001",
            "0000000000000001100001011001001111111111",
            "0000000000000000000000110100000010000011",
            "0000000000000001100000111000100001011111",
            "0000000000000001100001010000110001000001",
            "0000000000000001100001011001001111111111",
            "0000000000000001100000110001000010000011",
            "0000000000000000000000111100000010011111",
            "0000001100011101000000000111111111111111",
            "0000000000000001100000111000010000111111",
            "0000001100100101000000000111111111111111",
            "0000001100111110100000000000101111110000",
            "0000000000000001101000000111111111100001",
            "0000001000101001000000000100001111100101",
            "0000000000000001100100011111110010000010",
            "0000001010001101000000000111111111111111",
            "0000000000000010000000111100001111110000",
            "0000000000000001111000000111111111100010",
            "0000001101000111000000101001000010000100",
            "0000000000000001100000111000100001011111",
            "0000000000000001100000010001001111100100",
            "0000000000000001100000000100001111100100",
            "0000000000000001111000000100001111100011",
            "0000001101010001000000000111111111111111",
            "0000000000000001100000111000110001111111",
            "0000000000000001100000010001001111100100",
            "0000000000000011100000000000011111111111",
            "0000000000000001100000000001011111111111",
            "0000000000000001100100110000110001100011",
            "0000001101110111001100111111110001000011",
            "0000001101010101000000110000010000100001",
            "0000000000000001101100111111110001100010",
            "0000001101100011000000000111111111111111",
            "0000000000000001100000111000100001100010",
            "0000000000000001100000110001010000100101",
            "0000000000000001110011000000011111100001",
            "0000001101011011000011000000111111100011",
            "0000000000000001100100000111111111100100",
            "0000001101101101000000000111111111111111",
            "0000000000000001100000111001010010111111",
            "0000000000000001100000000000111111110000",
            "0000000000000001100100000111111111110000",
            "0000001101110101000000000111111111111111",
            "0000000000000001100000111000100001011111",
            "0000000000000000000000000000011111111111",
            "0000000000000001100000000000111111110000",
            "0000000000000001100000000001001111110000",
            "0000000010000010000000000000011111111111",
            "0000001110100111000100000000011111110000",
            "0000001110100111011000000111111111100010",
            "0000001110001111000000000111111111111111",
            "0000000001000001101100110111111111100010",
            "0000001110001001000011110000010001000001",
            "0000000000000000000000000100001111111111",
            "0000000000000011100011110000110001011111",
            "0000000000000011100000111000111111100011",
            "0000000000000000000001000100000001100001",
            "0000000001000001101100111111111111100010",
            "0000001110010111011000000111111111100001",
            "0000001110100111000000101000010000100001",
            "0000000000000000000000010100001111100001",
            "0000001110100001000011110000010001000001",
            "0000000000000011100011110000110001011111",
            "0000000000000011100000111000111111100011",
            "0000000000000001100000010000111111100011",
            "0000000000000000000000100100000001100001",
            "0000000000000011100011110000110001011111",
            "0000000000000011100000111000111111100011",
            "0000000000000000000000011100000001100001",
            "0000000000000000000000000100001111100001",
            "0000000000000001100000110000011000010100",
            "0000000000000000000010000100001010100001",
            "0000000000000001100000000000101111110000",
            "0000000000000001100000110000011000010100",
            "0000000000000000000010000101100001000001",
            "0000000000000011100011111000101111110000",
            "0000000000000011100011111000011111110000",
            "0000000000000011100000000001111111111111",
            "0000000000000111100001110111111111111111",
            "0000000000000001101011010000111111100001",
            "0000001111000011000000000111111111111111",
            "0000000000000001100000000001111111111111",
            "0000000000000011100000000000111111111111",
            "0000000000000001100010000000010011100001",
            "0000000000000011100000011001011111100001",
            "0000000000000011100001000000011111100001",
            "0000000000000001100000110000010000100001",
            "0000000000000011100000000001111111111111",
            "0000000000000111100001110111111111111111",
            "0000000000000001101011010001001111100010",
            "0000001111010111000000000111111111111111",
            "0000000000000001100000000001111111111111",
            "0000000000000011100000000001001111111111",
            "0000000000000001100010000000100011100010",
            "0000000000000011100000011001101111100010",
            "0000000000000011100001000000101111100010",
            "0000000000000000000000110000100001000010",
            "0000000000000001100000000000011111111111",
            "0000000000000001101000000111111111100001",
            "0000001111101011000000000111111111111111",
            "0000000000000001100000100000010010100001",
            "0000000000000011100011110000011111100001",
            "0000000000000000000000000100001111100001",
            "0000000000000001100000000001111111111111",
            "0000000000000111100001110111111111100111",
            "0000000000000101100010000001111111100111",
            "0000000000000001100000110010000011100111",
            "0000000000000001101100111111110100000001",
            "0000001111111011000000000111111111111111",
            "0000000000000011100000110000111111100011",
            "0000001111110011000011011000011111100001",
            "0000000000000001111000000111111111100011",
            "0000010000000011000000000111111111111111",
            "0000000000000011100000110000111111100011",
            "0000001111111011000011011000011111100001",
            "0000000000000001101000000111111111100011",
            "0000010000001011000000000111111111111111",
            "0000000000000011100000110000111111100011",
            "0000000000000001100011011000011111100001",
            "0000000000000001110000111111110011100001",
            "0000010000010111000000000111111111111111",
            "0000000000000011100100111111111111100011",
            "0000010000010111000000000111111111111111",
            "0000000000000011100000111000111111100011",
            "0000010000001011000000110000010000100001",
            "0000000000001001100100011111111111100001",
            "0000010000011101000000000111111111111111",
            "0000000000000011100000110000011111100001",
            "0000000000000011100000110000011111100001",
            "0000000000000001101100111111110100000001",
            "0000010000100111000000000111111111111111",
            "0000000000000011100000110000111111100011",
            "0000010000010111000011011000011111100001",
            "0000000111111111110000111111111111100011",
            "0000010001000101010000111111110011100001",
            "0000010000101111000000000111111111111111",
            "0000000000000001100000000000111111111111",
            "0000000000000001100011000000011111100001",
            "0000000000000011100101000000011111100001",
            "0000010001010001000000000111111111111111",
            "0000000000000111100001110111111111111111",
            "0000001111100101000010000000010001100001",
            "0000000000000001100010111000011111111111",
            "0000000000000001100010000000011111100001",
            "0000000110000001100010000000011111100001",
            "0000000111111111100010000100001111100001",
            "0000000010000101100000000000011111111111",
            "0000001000101001000000000111111111111111",
            "0000000000000111100001110111111111111111",
            "0000000111111111100010000000011111100101",
            "0000000000000011100011110000011111100001",
            "0000000000000001100000000100001111100001",
            "0000000010000101100000000000011111111111",
            "0000001000101001000000000111111111111111",
            "0000000000000011100011110100001111100101",
            "0000000010000111100000000000011111111111",
            "0000001000101001000000000111111111111111",
            "0000010100101100100000000111111111111111",
            "0000001110110010100000000111111111111111",
            "0000000000000001100100000111111111100010",
            "0000010010001111010000111001110010000011",
            "0000010001110001000000111010000001100100",
            "0000000000110101101100111111111111101000",
            "0000010001101011000000000111111111111111",
            "0000000000000001100000000000011111100010",
            "0000000000000001100000000000111111100100",
            "0000001111100001000000000001011111100110",
            "0000000000000011101000111010001111101000",
            "0000010001101011000011000000011111100001",
            "0000010001111011000000000000111111100100",
            "0000000000110101110000111111111111100111",
            "0000001111100001000100000111111111100111",
            "0000010001111011000000000111111111111111",
            "0000000000000011101000111001111111100111",
            "0000010001110111000011000000101111100010",
            "0000000000000001100100000111111111100101",
            "0000010010000001000000000111111111111111",
            "0000000000000001100000111000010000111111",
            "0000000000000001100100000111111111100110",
            "0000010010000111000000000111111111111111",
            "0000000000000001100000111000100001011111",
            "0000000000000001111000110000010001000001",
            "0000001111100001000010110001010010100101",
            "0000000000000001100000111000010000111111",
            "0000001111100001000010101001010010100101",
            "0000000000000001101000000111111111100001",
            "0000001111100001000000000111111111111111",
            "0000001111100001000000011001010011000101",
            "0000001110110010100000000111111111111111",
            "0000000000000001100000101001010011000101",
            "0000000000000001100100000111111111100001",
            "0000001111100001000100000111111111100010",
            "0000001111011111000000000111111111111111",
            "0000000000000001100000110000110010000011",
            "0000000100110001100000111000111111100011",
            "0000000000000001100000000010001111111111",
            "0000000000000111100001110111111111101000",
            "0000000000000101100010000010001111101000",
            "0000000000000001100000000001111111100001",
            "0000000000000001100000000000011111111111",
            "0000000000000001110011000000101111100010",
            "0000010010110011000000000111111111111111",
            "0000000000000001100000110000010011100001",
            "0000000000000001100100000111111111100010",
            "0000001111100001010000111111110100000111",
            "0000010010111011000000000111111111111111",
            "0000010010101101000000110001110011100111",
            "0000000000000011100000110000111111100011",
            "0000010010101101000011000000011111100001",
            "0000001110110010100000000111111111111111",
            "0000000000000001100000101001010011000101",
            "0000000000000001100100000111111111100010",
            "0000010011111011000100000111111111100001",
            "0000001111100001000000000111111111111111",
            "0000000000000001100000111000110010000011",
            "0000000011111011100000110000111111100011",
            "0000000000000001100000000010001111111111",
            "0000000000000111100001110111111111101000",
            "0000000000000101100010000010001111101000",
            "0000000000000001110000111111110100000001",
            "0000010011011011000000000111111111111111",
            "0000000000000011100000111000111111100011",
            "0000010011010011000000110000010000100001",
            "0000000000000001110000111111110100000010",
            "0000010011100011000000000111111111111111",
            "0000000000000011100000110000111111100011",
            "0000010011011011000000110000100001000010",
            "0000000000000001100000000001111111100001",
            "0000000000000001100000000000011111111111",
            "0000000000111001100000000010001111111111",
            "0000000000000001101100111111110001000111",
            "0000010011110001000000110000010000100001",
            "0000000000000001100000111001110001000111",
            "0000000000000011100000110000011111100001",
            "0000000000000011101000111010001111101000",
            "0000010011101001000100110001110011100111",
            "0000001111100001000000000111111111111111",
            "0000000000000011100000100000011111100001",
            "0000001111100001000000000111111111111111",
            "0000010000111001000000000111111111111111",
            "0000010001000101000000000111111111111111",
            "0000000000000001100000000000101111110000",
            "0000000000000001100000000000011111110000",
            "0000000000000011100011110000111111111111",
            "0000000000000001100001000001010001100001",
            "0000000000000001100001000001100001100010",
            "0000000000000001100010100000110011000101",
            "0000000000000001100010010001000011000101",
            "0000000000000001101000000111111111100101",
            "0000010100010011000000000111111111111111",
            "0000000000000001100000000000111111111111",
            "0000000000000001101000000111111111100110",
            "0000010100011001000000000111111111111111",
            "0000000000000001100000000001001111111111",
            "0000000000000001111000000111111111100001",
            "0000010100011111000000000111111111111111",
            "0000000000000001100000111000110001111111",
            "0000000000000001111000000111111111100010",
            "0000010100100101000000000111111111111111",
            "0000000000000001100000111001000010011111",
            "0000000000000001100000000100001111100011",
            "0000000000000000000000000100001111100100",
            "0000000000000011100011110000011111111111",
            "0000000000000000000001000100000000110000",
            "0000000000000011100011110000011111111111",
            "0000000000000000000000101100000000110000",
            "0000000000000001100100001000011001111111",
            "0000010100111101000000000111111111111111",
            "0000000000000011100100111111111111100001",
            "0000010101001001000000000111111111111111",
            "0000000000000101100000111100101111110010",
            "0000001000010001000000000111111111111111",
            "0000000000000001100000000000011111110000",
            "0000000100110001100000000000111111111111",
            "0000000000000001111000000111111111100001",
            "0000001111100001000010110001010010100101",
            "0000000000000001100000111000010000111111",
            "0000001111100001000010101001010010100101",
            "0000000000000011100011111000101111110000",
            "0000001111001010100000000111111111111111",
            "0000000011111111110000111111111111100100",
            "0000010101010101000000000111111111111111",
            "0000000000000001100000000000101111111111",
            "0000000000000000000000000100001111100010",
            "0000000100110001110000111111111111100100",
            "0000010101011101000000000111111111111111",
            "0000000000000011100000110001001111100100",
            "0000010101010101000011000000101111100010",
            "0000000100110001100100111111111111100100",
            "0000010101101011000000000111111111111111",
            "0000000000000011100000111001001111100100",
            "0000000000000001111000110000100001000010",
            "0000010101011101000000000111111111111111",
            "0000000000000011100011110000101111100110",
            "0000001000010101000000000100001111100010",
            "0000000000000001100100000111111111100110",
            "0000010101010011000000000111111111111111",
            "0000000000000001100000111000100001011111",
            "0000010101010011000000000111111111111111",
            "0000010101110111000000000111111111111111",
            "0000000000000000000000111100000000111111",
            "0000000000000000000000000100001111100001",
            "0000000000000001100000000000101111110000",
            "0000000000000011100011111000010001011111",
            "0000000001000001110000111111111111100010",
            "0000010110000011000000011000010001100001",
            "0000000000000000000010110100000000111111",
            "0000000000000000000000000100001111111111",
            "0000000001000001110000111111111111100010",
            "0000001000011111000000000111111111111111",
            "0000000000000010000011111100000001011111",
            "0000001100111110100000000000101111110000",
            "0000000000000001101000000111111111100001",
            "0000001000101001000000000100001111100010",
            "0000000000000001100100011111110010000010",
            "0000001010001101000000000111111111111111",
            "0000000000000000000000110100000001110000",
            "0000000111011000100000000001011111110000",
            "0000000000000000000000000100001111100101",
            "0000000110110100100000000001011111110000",
            "0000000000000001100000000101100010101110",
            "0000000000000010000000110011101111101110",
            "0000000000000001100011000000011111110000",
            "0000000000000001100011000100001111100001",
            "0000000000000011100000110000011111110000",
            "0000000000000001100000110000101001101100",
            "0000000000000001100000000101100111000010",
            "0000000000000001100000000000101111110000",
            "0000000000000001100000000000111010100010",
            "0000000000000001100000000101100001101110",
            "0000000000000011100000110011101111101110",
            "0000000000000011100000110000101111100010",
            "0000000000000011101000111000011111100001",
            "0000010110101101000000000111111111111111",
            "0000000000000000000000000111111111111111",
            "0000000000000001100010111000011001111111",
            "0000000000000001100010000000011001100001",
            "0000000000000001100000110100100000110010",
            "0000001010001100100000000000011111110000",
            "0000000000000001100010111000101001111111",
            "0000000000000001100010000000101001100010",
            "0000000000000001100010111000111001111111",
            "0000000000000001100010000000111001100011",
            "0000000000000001100000111001000001000011",
            "0000000000000001100000110001000010000100",
            "0000000000001001100000110001001111100100",
            "0000000000000001100000110001001001000100",
            "0000000000000001100000000101100010001110",
            "0000000000000011100000110011101111101110",
            "0000000000000001100010100001000001000001",
            "0000000000000001100010010001010001100001",
            "0000000000000001100100011111110010100100",
            "0000010111100101000000111000010001000001",
            "0000000000000011100000110000011111100001",
            "0000000000000001100000110000010000100001",
            "0000001010001010100000110100100000110010",
            "0000000000000001100010111000011001111111",
            "0000000000000001100010000000011001100001",
            "0000001010001001000000111100100000110010",
            "0000000000000011100000111011101111101110",
            "0000000000000001100000000100101010101110",
            "0000001010001011000000000111111111111111",
            "0000000000000001100010000000011001100001",
            "0000000000000001100000110000010000110010",
            "0000000000000001100000000101100000101110",
            "0000000000000010000000110011101111101110",
            "0000111000110111000000000111111111111111",
            "0000001010001101000000000111111001110000",
            "0000000000000001100000000000101111110000",
            "0000000000000111100100011001001111100011",
            "0000011000001111000000000000011111110000",
            "0000000000000001100000000001011010100010",
            "0000000000000001100000000101100010100001",
            "0000000000000011100000110000011111100001",
            "0000000000000011100000110000101111100010",
            "0000000000000011101000111001001111100100",
            "0000011000000011000000000111111111111111",
            "0000000000000111100101000001001111100011",
            "0000001010001101000000000111111111111111",
            "0000000000000001100000000001011010100010",
            "0000000000000001100000000101100010100001",
            "0000000000000001100000001001011010100010",
            "0000000000000001100000001101100010100001",
            "0000000000000001100000010001011010100010",
            "0000000000000001100000010101100010100001",
            "0000000000000001100000011001011010100010",
            "0000000000000001100000011101100010100001",
            "0000000000001001100000110000011111100001",
            "0000000000001001100000110000101111100010",
            "0000000000001001101000111001001111100100",
            "0000011000010011000000000111111111111111",
            "0000000000000000000000000111111111111111",
            "0000000000000001110000111111111101100001",
            "0000001000001101000000000100001111100001",
            "0000000000000000000000000111111111111111",
            "0000000000000001100010000000101001100010",
            "0000000000000001100000001000011010101011",
            "0000000000000000000000110100000001000001",
            "0000000000000001100001110000011111110000",
            "0000000000000001100000000100001111100110",
            "0000000000000001100000000001011010100001",
            "0000000000000001100000000001101010100010",
            "0000000000000011100000110000011111100001",
            "0000000000000011100000110000101111100010",
            "0000000000000001100111010000111111100101",
            "0000011001100101000001111001001111100110",
            "0000000000000001101000101111110010000011",
            "0000011001100101000000000111111111111111",
            "0000000000000001100111010000111111100101",
            "0000011001100101000001111001001111100110",
            "0000000000000001101000101111110010000011",
            "0000011001100101000000000111111111111111",
            "0000000000000001100111010000111111100101",
            "0000011001100101000001111001001111100110",
            "0000000000000001101000101111110010000011",
            "0000011001100101000000000111111111111111",
            "0000000000000001100111010000111111100101",
            "0000011001100101000001111001001111100110",
            "0000000000000001100100101111110010000011",
            "0000011000111101000000000111111111111111",
            "0000000000000001100000000001101111110000",
            "0000000000000001100000000100001111100011",
            "0000000000000000000000000100001111100100",
            "0000000000000001100000000000011111101100",
            "0000000000000001100100001000101001111111",
            "0000011001110111000000000111111111111111",
            "0000000000000001100000000000011010100001",
            "0000000000000011101000111000101111100010",
            "0000011001110001000000000111111111111111",
            "0000000000000000000000000100001111100001",
            "0000000000000001100000000000101111110000",
            "0000000000000001100000000000011111110000",
            "0000000000000001100010100001000001000001",
            "0000000000000001100010010001010001100001",
            "0000000000000001100100011111110010100100",
            "0000001000100001000000000100001111100001",
            "0000000000000000000000000111111111111111",
            "0000000000000001100000000000011111110000",
            "0000000000000001100010100001001111100001",
            "0000000000000001100010010001010001000001",
            "0000000000000001100100011111110010100100",
            "0000001000100001000000000100001111100001",
            "0000000000000000000000000111111111111111",
            "0000000000000001100000000100001111101110",
            "0000000000000000000000110011100000101110",
            "0000000000000001111000000111111111100001",
            "0000011010011111000000000011101111101100",
            "0000000000000001100000000010111010101110",
            "0000000000000001100000000011111010101011",
            "0000000000000001100000000100101111100001",
            "0000000000000001100000001011001010101110",
            "0000001010001101000000000111111111111111",
            "0000000000000001100000111000011001101011",
            "0000000000000011100000111000011111100001",
            "0000000000000001100000000000011010100001",
            "0000000000000001100000001000101001111111",
            "0000000000000011100011110000111111111111",
            "0000000000000001100000100000110001110010",
            "0000000000000001100000000101100101101110",
            "0000000000000001100000001101100110001110",
            "0000000000000001100000010101100001101110",
            "0000000000000001100000000011001111101110",
            "0000000000001001100000110011101111101110",
            "0000000000000001100000000010111010100001",
            "0000000000000001100000000011111010101011",
            "0000000000000001100000110000100001001111",
            "0000000000000001100000000100101010100010",
            "0000001010001011000000000111111111111111",
            "0000000000000001100000110000011001101111",
            "0000000000000001100000000101101000001110",
            "0000011011011001000000000111111111111111",
            "0000000000000011100000111011101111101110",
            "0000000000000001100000000000011010101110",
            "0000000000000001100000000000111111111111",
            "0000000000000111100001110111111111100011",
            "0000000000000001100011010000101111100001",
            "0000011010101101000010000000010001100001",
            "0000000000000001100000000101100110001110",
            "0000000000000001100000010101101001001110",
            "0000000000000001100000000100101010100001",
            "0000000000000001100000001101100110001110",
            "0000000000000001100000000011001111101110",
            "0000000000001000000000110011101111101110",
            "0000000001000001110000111111111111100010",
            "0000001000011101000000000000111111110000",
            "0000000000000011100011111000010001011111",
            "0000000000000001100000000001001010100011",
            "0000000000000001100000100001000000100100",
            "0000000000000000000000000101100010000011",
            "0000000001000001110000111111111111100010",
            "0000001000011101000000000000111111110000",
            "0000000000000011100011111000010001011111",
            "0000000000000001100000000001001010100011",
            "0000000000000001100001000001000000100100",
            "0000000000000000000000000101100010000011",
            "0000000000000001100000000000101111110000",
            "0000000000000001100000000000011111110000",
            "0000000000000001111000111111110001100001",
            "0000011100000101000000000111111111111111",
            "0000000000000000000000000100001111111111",
            "0000000000000011100011111000110000111111",
            "0000000000111111100001000000011111100001",
            "0000000000001011100011110000011111100001",
            "0000000000000001100000110000010000100010",
            "0000000000000001100000000001001010100001",
            "0000000000000001100000011000110010000011",
            "0000000000000000000010110100001111100011",
            "0000000000000001100000000000101111110000",
            "0000000000000011100000000001001111111111",
            "0000000000000001100100001000011001111111",
            "0000011100100111000100111000010010000001",
            "0000011100101001000100111000010010000001",
            "0000011100110001000100111000010010000001",
            "0000011100110011000000000111111111111111",
            "0000000000000001100000000100001111100010",
            "0000000000000001100000000100001111100011",
            "0000001000010001000000111100100010010010",
            "0000001000010001000000000111111111111111",
            "0000001100111110100000000111111111111111",
            "0000000000000001101000000111111111100001",
            "0000001000101001000000000100001111100101",
            "0000000000000000000000000111111111111111",
            "0000001000010001000000000111111111111111",
            "0000001100111110100000000111111111111111",
            "0000000000000001101000000111111111100001",
            "0000001000101001000000000100001111100010",
            "0000000000000000000000000111111111111111",
            "0000000000000001100000000000101010100001",
            "0000000000000011100000110000101111100010",
            "0000000000000000000000000101100001000001",
            "0000000000000001100000000000101010100001",
            "0000000000000011100000111000101111100010",
            "0000000000000000000000000101100001000001",
            "0000000000000001100000000000011111110000",
            "0000000000000001100000000000111010100001",
            "0000000000000001100000110000110001000011",
            "0000000000000000000000000101100001100001",
            "0000000000000001100000000000011111110000",
            "0000000000000001100000000000111010100001",
            "0000000000000001100000111000110001000011",
            "0000000000000000000000000101100001100001",
            "0000000000000001100000000101101000001110",
            "0000000000000010000000110011101111101110",
            "0000000000000011100000111011101111101110",
            "0000000000000000000000000100001010101110",
            "0000000000000001100001011000101111111111",
            "0000000000000001100000110000100001000001",
            "0000000000000000000000110100000001010000",
            "0000000000000001100000001000101001111111",
            "0000000000000001100000111000010000101011",
            "0000000000000011100000111000011111100001",
            "0000000000000001100000000000011010100001",
            "0000000000000111100001110111111111111111",
            "0000000000000000000010000100000001000001",
            "0000000000000001100000000000011111110000",
            "0000000000000001100000000000111010100001",
            "0000000000000001100000001001001010100001",
            "0000000000000001100000000100001111100011",
            "0000000000000001100000000100001111100010",
            "0000000000000001100010011001000010000010",
            "0000000000000001100010001001011111100010",
            "0000000000000001100100100111110010100100",
            "0000001010001101000000000111111111111111",
            "0000001000100001000000000111111111111111",
            "0000000000000000000000000100001111111100",
            "0000000000000010000000111100001111100001",
            "0000000000000011100000111000011111100001",
            "0000000000000000000000000100001010100001",
            "0000000000000011100000111000011111100001",
            "0000000000000000000000000101101000000001",
            "0000000000000001100000000000011111110000",
            "0000000000000001100000000101100001000001",
            "0000000000000000000000000100001111100010",
            "0000000000000001100000000000101111110000",
            "0000000000000001100000000000011111110000",
            "0000000000000001100010100001000001000001",
            "0000000000000001100010010001010001100001",
            "0000000000000000000000011100000010100100",
            "0000000000000001100000000000011111110000",
            "0000000000000001100010100001001111100001",
            "0000000000000001100010010001010001000001",
            "0000000000000000000000011100000010100100",
            "0000000000000011100000111011101111101110",
            "0000000000000001100000000000011010101110",
            "0000000000000011100011110000111111111111",
            "0000000000000001100000100000110001110010",
            "0000000000000001100000000101100101101110",
            "0000000000000001100000001101100110001110",
            "0000000000000001100000010101100001101110",
            "0000000000000001100000000011001111101110",
            "0000000000001001100000110011101111101110",
            "0000011010111101000000000010111111100001",
            "0000000000000001100000001000011001111111",
            "0000000000000001100100111111111111100001",
            "0000011111001111000000000111111111111111",
            "0000000000000011100100111111111111100001",
            "0000011111010001000000000111111111111111",
            "0000000000000101100100111111111111100001",
            "0000011111011001000000000111111111111111",
            "0000000000000011100000111100101111110010",
            "0000001000010001000000000111111111111111",
            "0000000000001110000000000100001111111111",
            "0000000000000001100000000000011111110000",
            "0000000110010000100000000111111111111111",
            "0000000000011011100000000101101111110100",
            "0000000000010100000000000101101111110100",
            "0000000000000000000000000100001111111111",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000000000000000000000000000000000",
            "0000000000100001100000000000011111111111",
            "0000001001011111000000000111111111111111",
            "0000000000000011100000000000011111111111",
            "0000001001011111000000000111111111111111",
            "0000000000100101100000000000011111111111",
            "0000001001011111000000000111111111111111",
            "0000000000100111100000000000011111111111",
            "0000001001011111000000000111111111111111",
            "0000000000101001100000000000011111111111",
            "0000001001011111000000000111111111111111",
            "0000000000101011100000000000011111111111",
            "0000001001011111000000000111111111111111",
            "0000000000101101100000000000011111111111",
            "0000001001011111000000000111111111111111",
            "0000000000101111100000000000011111111111",
            "0000001001011111000000000111111111111111",
            "0000001001100101000000000111111111111111",
            "0000001010000011000000000111111111111111",
            "0000001010000101000000000111111111111111",
            "0000001010000101000000000111111111111111",
            "0000001010000101000000000111111111111111",
            "0000001010000101000000000111111111111111",
            "0000001010000101000000000111111111111111",
            "0000001010000101000000000111111111111111",
            "0000001010000101000000000111111111111111",
            "0000001010000101000000000111111111111111",
            "0000001010000101000000000111111111111111",
            "0000001010000101000000000111111111111111",
            "0000001010000101000000000111111111111111",
            "0000001010000101000000000111111111111111",
            "0000001010000101000000000111111111111111",
            "0000001010000101000000000111111111111111",
            "0000000000000000000000000100001111111111",
            "0000000000000010000000000100001111111111",
            "0000000000000100000000000100001111111111",
            "0000000000000110000000000100001111111111",
            "0000000000001000000000000100001111111111",
            "0000000000001010000000000100001111111111",
            "0000000000001100000000000100001111111111",
            "0000000000001110000000000100001111111111",
            "0000000000010000000000000100001111111111",
            "0000000000010010000000000100001111111111",
            "0000000000010100000000000100001111111111",
            "0000000000010110000000000100001111111111",
            "0000000000011000000000000100001111111111",
            "0000000000011010000000000100001111111111",
            "0000000000011100000000000100001111111111",
            "0000000000011110000000000100001111111111",
            "0000001010001101000000001100001001111111",
            "0000001010001111000010111000011001111111",
            "0000001010010001000010111000011001111111",
            "0000000000000000000000001100001101111111",
            "0000001010001101000000110100001001101100",
            "0000001010001101000000110100001001101011",
            "0000001010001101000000110100001001110000",
            "0000001010010111000000111000011001101011",
            "0000001010100001000100000111111111110000",
            "0000001010100101000000000111111111111111",
            "0000001010101011000100000111111111110000",
            "0000001010001011000000000111111111111111",
            "0000001010101111000100000111111111110000",
            "0000001010110011000000000111111111111111",
            "0000001010111001000100000111111111110000",
            "0000001010001011000000000111111111111111",
            "0000001010111101000000110000011001101100",
            "0000001010111111000000110000011001101011",
            "0000001011000001000000111000011001101011",
            "0000001011001011000000110000011001110000",
            "0000000000000000000000100100001010101100",
            "0000000000000000000000101100001010101100",
            "0000000000000000000000110100001010101100",
            "0000000000000000000000111100001010101100",
            "0000000000000000000001000100001010101100",
            "0000000000000000000001001100001010101100",
            "0000000000000000000001010100001010101100",
            "0000000000000000000001011100001010101100",
            "0000000000000000000001100100001010101100",
            "0000000000000000000001101100001010101100",
            "0000000000000000000001110100001010101100",
            "0000000000000000000001111100001010101100",
            "0000001011001101000000110000011001101100",
            "0000001011001111000000110000011001101011",
            "0000001011010001000000111000011001101011",
            "0000001011011011000000000000101111110000",
            "0000000000000000000000100101101000001100",
            "0000000000000000000000101101101000001100",
            "0000000000000000000000110101101000001100",
            "0000000000000000000000111101101000001100",
            "0000000000000000000001000101101000001100",
            "0000000000000000000001001101101000001100",
            "0000000000000000000001010101101000001100",
            "0000000000000000000001011101101000001100",
            "0000000000000000000001100101101000001100",
            "0000000000000000000001101101101000001100",
            "0000000000000000000001110101101000001100",
            "0000000000000000000001111101101000001100",
            "0000001011011111000001110000011000010000",
            "0000001011100011000000110000011000010000",
            "0000000000000000000000010100001010101011",
            "0000000000000000000000011100001010101011",
            "0000000000000000000000100100001010101011",
            "0000000000000000000000101100001010101011",
            "0000000000000000000000110100001010101011",
            "0000000000000000000000111100001010101011",
            "0000000000000000000001000100001010101011",
            "0000000000000000000001001100001010101011",
            "0000000000000000000001010100001010101011",
            "0000000000000000000001011100001010101011",
            "0000000000000000000001100100001010101011",
            "0000000000000000000001101100001010101011",
            "0000000000000000000001110100001010101011",
            "0000000000000000000001111100001010101011",
            "0000001011100101000000000000111111110000",
            "0000001011101101000000000000101111110000",
            "0000000000000000000000010101101000001011",
            "0000000000000000000000011101101000001011",
            "0000000000000000000000100101101000001011",
            "0000000000000000000000101101101000001011",
            "0000000000000000000000110101101000001011",
            "0000000000000000000000111101101000001011",
            "0000000000000000000001000101101000001011",
            "0000000000000000000001001101101000001011",
            "0000000000000000000001010101101000001011",
            "0000000000000000000001011101101000001011",
            "0000000000000000000001100101101000001011",
            "0000000000000000000001101101101000001011",
            "0000000000000000000001110101101000001011",
            "0000000000000000000001111101101000001011",
            "0000000000000000000000000100001010110000",
            "0000000000000000000000001100001010110000",
            "0000000000000000000000010100001010110000",
            "0000000000000000000000011100001010110000",
            "0000000000000000000000100100001010110000",
            "0000000000000000000000101100001010110000",
            "0000000000000000000000110100001010110000",
            "0000000000000000000000111100001010110000",
            "0000000000000000000001000100001010110000",
            "0000000000000000000001001100001010110000",
            "0000000000000000000001010100001010110000",
            "0000000000000000000001011100001010110000",
            "0000000000000000000001100100001010110000",
            "0000000000000000000001101100001010110000",
            "0000000000000000000001110100001010110000",
            "0000000000000000000001111100001010110000",
            "0000000000000000000000000101101000010000",
            "0000000000000000000000001101101000010000",
            "0000000000000000000000010101101000010000",
            "0000000000000000000000011101101000010000",
            "0000000000000000000000100101101000010000",
            "0000000000000000000000101101101000010000",
            "0000000000000000000000110101101000010000",
            "0000000000000000000000111101101000010000",
            "0000000000000000000001000101101000010000",
            "0000000000000000000001001101101000010000",
            "0000000000000000000001010101101000010000",
            "0000000000000000000001011101101000010000",
            "0000000000000000000001100101101000010000",
            "0000000000000000000001101101101000010000",
            "0000000000000000000001110101101000010000",
            "0000000000000000000001111101101000010000",
            "0000000000000000000000000111111111111111",
            "0000000000101001000000000111111111111111",
            "0000000000000000000000000100001111101101",
            "0000001011110001000000000011011111110000",
            "0000001000101001000000000000011111110000",
            "0000001011111101000000000001011111110000",
            "0000001100001101000000000000011111110000",
            "0000001100010001000000000111111111111111",
            "0000000000000000000000110100001000010000",
            "0000000000000000000000111100001000010000",
            "0000001100010101011000000000101111110000",
            "0000001100110011000000000000111111110000",
            "0000000000000001100000111100001000011111",
            "0000001101111101000100000000101111110000",
            "0000000000000000000011111100001000010000",
            "0000000000000000000011110100001000010000",
            "0000001000010001000000000111111111111111",
            "0000001000010001000000000111111111111111",
            "0000000000000000000000000100001010110100",
            "0000000000000000000000000101101000010100",
            "0000001000010001000000000111111111111111",
            "0000001000010001000000000111111111111111",
            "0000001110101001000000000111111111111111",
            "0000001110101101000000000111111111111111",
            "0000010001011001000000000111111111111111",
            "0000010001010111000000000111111111111111",
            "0000010010010101000000000111111111111111",
            "0000010010111111000000000111111111111111",
            "0000010011111111000000000111111111111111",
            "0000010100101001000000000111111111111111",
            "0000010100101101000000000111111111111111",
            "0000010100110001000000000111111111111111",
            "0000000000000000000010001100001000010000",
            "0000000000000000000010010100001000010000",
            "0000000000000000000010011100001000010000",
            "0000000000000000000010100100001000010000",
            "0000000000000000000010101100001000010000",
            "0000000000000000000010110100001000010000",
            "0000010101110011011000000000011111110000",
            "0000000000000000000000111100001000011111",
            "0000000000000000000000100100001000010000",
            "0000000000000000000000011100001000010000",
            "0000000000000000000000101100001000010000",
            "0000000000000000000001000100001000010000",
            "0000010101111001000000000000111111110000",
            "0000010110000101000000000000101111110000",
            "0000000000000000000010101100001111110000",
            "0000010110001011000000000000111111110000",
            "0000000000000000000000111011101000001110",
            "0000000000000000000000000111111111110000",
            "0000010110010111000000000111111111111111",
            "0000000110110101000000000111111111111111",
            "0000010110011011000000000111111111111111",
            "0000000000000000000000000100001101010000",
            "0000010110100001000000000111111111111111",
            "0000010110100101000000000111111111111111",
            "0000001000010001000000000111111111111111",
            "0000001000010001000000000111111111111111",
            "0000010110111011000000000111111111111111",
            "0000010111101011000000000111111111111111",
            "0000010111110001000010111000011001111111",
            "0000001010001001000000000100101111110000",
            "0000010111111001001000000100001111110000",
            "0000010111111001000100000100001111110000",
            "0000010111111101000000000000111111110000",
            "0000011000101101000000000000011111110000",
            "0000011000110011000010111000101001111111",
            "0000011000111001000000000000101111110000",
            "0000011001101011000000000111111111111111",
            "0000000000000000000000000100001010101100",
            "0000011001111001000000000000111111110000",
            "0000011010000111000000000000101111110000",
            "0000011010010011000000000000011111110000",
            "0000001010001101000000110011101001101110",
            "0000011010010111000000010000011010101100",
            "0000000000000000000000000111111111111111",
            "0000011010100101000000000111111111111111",
            "0000011011000101000000000111111111111111",
            "0000011011001011000000000111111111111111",
            "0000011011010111000000110000011001101111",
            "0000011011010111000000110000010111110011",
            "0000011011010111000000110000010111110011",
            "0000011011010111000000110000010111110011",
            "0000011011010111000000110000010111110011",
            "0000011011010111000000110000010111110011",
            "0000011011010111000000110000010111110011",
            "0000011011010111000000110000010111110011",
            "0000011011010111000000110000010111110011",
            "0000011011010111000000110000010111110011",
            "0000011011010111000000110000010111110011",
            "0000011011010111000000110000010111110011",
            "0000011011010111000000110000010111110011",
            "0000011011010111000000110000010111110011",
            "0000011011010111000000110000010111110011",
            "0000011011010111000000110000010111110011",
            "0000011011010111000000110000010111110011",
            "0000011011100011000000000000101111110000",
            "0000011011101111000000000000101111110000",
            "0000011011111011000000000000111111110000",
            "0000011100010011000000000000111111110000",
            "0000011100111011000000000000011111110000",
            "0000011101000001000000000000011111110000",
            "0000011101000111000000000000101111110000",
            "0000011101001111000000000000101111110000",
            "0000011101010111000000000111111111111111",
            "0000011101011011000000000111111111111111",
            "0000011101011111000001010000011000010000",
            "0000011101100101000000001000011001111111",
            "0000001000010001000000000111111111111111",
            "0000001000010001000000000111111111111111",
            "0000001000010001000000000111111111111111",
            "0000011101110001000000000000101111110000",
            "0000011110000101000000001100001000010000",
            "0000011110000111000000111000011001101100",
            "0000011110001001000000111000011001101100",
            "0000011110001101000000111000011001101100",
            "0000011110010001000000000000101111110000",
            "0000011110010111000000000000111111110000",
            "0000011110100001000000000000101111110000",
            "0000011110101001000000001000101001111111",
            "0000001000010001000000000111111111111111",
            "0000001000010001000000000111111111111111",
            "0000000000000000000000000100001111101010",
            "0000001000010001000000000111111111111111",
            "0000011110111101000000000111111111111111",
            "0000001000010001000000000111111111111111",
            "0000011111010011000000000000011111110000",
            "0000001000011001000000000111111111111111"
            -- microcode end
            );
    begin
       	if clock'event and clock = '1' and en = '1' then
            data <= rom(conv_integer(addr));
 	end if;
    end process;

end Behavioral;
