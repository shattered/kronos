library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

library unisim;
use unisim.vcomponents.all;

-- Note: XST cannot infer block RAM with two writable ports

entity BlockRam is
    -- mode : read-first
    -- clock: rise
    -- write enable: high
    -- clock enable: high
    port (
	clock  : in std_logic;
	en0    : in std_logic;
	en1    : in std_logic;
	we0    : in std_logic;
	we1    : in std_logic;
	a0     : in std_logic_vector(8 downto 0);
	a1     : in std_logic_vector(8 downto 0);
	di0    : in std_logic_vector(31 downto 0);
	di1    : in std_logic_vector(31 downto 0);
	do0    : out std_logic_vector(31 downto 0);
	do1    : out std_logic_vector(31 downto 0));
end BlockRam;


architecture Behaviour of BlockRam is
    signal DOA   : std_logic_vector(31 downto 0);
    signal DOB   : std_logic_vector(31 downto 0);
    signal DOPA  : std_logic_vector(3 downto 0);
    signal DOPB  : std_logic_vector(3 downto 0);
    signal ADDRA : std_logic_vector(8 downto 0);
    signal ADDRB : std_logic_vector(8 downto 0);
    signal CLKA  : std_logic;
    signal CLKB  : std_logic;
    signal DIA   : std_logic_vector(31 downto 0);
    signal DIB   : std_logic_vector(31 downto 0);
    signal DIPA  : std_logic_vector(3 downto 0);
    signal DIPB  : std_logic_vector(3 downto 0);
    signal ENA   : std_logic;
    signal ENB   : std_logic;
    signal SSRA  : std_logic;
    signal SSRB  : std_logic;
    signal WEA   : std_logic;
    signal WEB   : std_logic;

begin
   -- RAMB16_S36_S36: Virtex-II/II-Pro, Spartan-3/3E 512 x 32 + 4 Parity bits Dual-Port RAM
   -- Xilinx  HDL Language Template version 7.1i

   RAMB16_S36_S36_inst : RAMB16_S36_S36
   generic map (
      INIT_A  => X"000000000",  --  Value of output RAM registers on Port A at startup
      INIT_B  => X"000000000",  --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"000000000", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"000000000", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL" 
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA   => DOA,     -- Port A 32-bit Data Output
      DOB   => DOB,     -- Port B 32-bit Data Output
      DOPA  => DOPA,    -- Port A 4-bit Parity Output
      DOPB  => DOPB,    -- Port B 4-bit Parity Output
      ADDRA => ADDRA,   -- Port A 9-bit Address Input
      ADDRB => ADDRB,   -- Port B 9-bit Address Input
      CLKA  => CLKA,    -- Port A Clock
      CLKB  => CLKB,    -- Port B Clock
      DIA   => DIA,     -- Port A 32-bit Data Input
      DIB   => DIB,     -- Port B 32-bit Data Input
      DIPA  => DIPA,    -- Port A 4-bit parity Input
      DIPB  => DIPB,    -- Port-B 4-bit parity Input
      ENA   => ENA,     -- Port A RAM Enable Input
      ENB   => ENB,     -- PortB RAM Enable Input
      SSRA  => SSRA,    -- Port A Synchronous Set/Reset Input
      SSRB  => SSRB,    -- Port B Synchronous Set/Reset Input
      WEA   => WEA,     -- Port A Write Enable Input
      WEB   => WEB      -- Port B Write Enable Input
   );

    do0 <= DOA;
    do1 <= DOB;
    ADDRA <= a0;
    ADDRB <= a1;
    CLKA <= clock;
    CLKB <= clock;
    DIA <= di0; 
    DIB <= di1;
    DIPA <= "0000";
    DIPB <= "0000";
    ENA <= en0;
    ENB <= en1;
    SSRA <= '0';
    SSRB <= '0';
    WEA <= we0;
    WEB <= we1;

end architecture Behaviour;
